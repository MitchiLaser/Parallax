* Analog Frontend

.include libs/analog_frontend.sub
* Instantiate like this:
* XAFEn IN OUT AnalogFrontend

* This is a list of all the parameters in use
* Amplitudes of the sine wave: 15, 5, 2, 0.5
* Resistor of the amplifier (multiplexer): ???
* Resistor of the Ref voltage generator (multiplexer): ???

* try out the analog frontend on a sinusodial input signal
Vsource Vsource 0 SIN(0 15 1000)
.param pamp=1G
.param pref=10k
XAFE1 Vsource VAFEout1 AnalogFrontend

.tran 100ns 2ms

.control
run
plot v(Vsource) v(VAFEout1) title "input and output voltage"
.endc
.end

